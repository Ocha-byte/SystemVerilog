`timescale 1 ns / 1ns

module alu (
    //input in1,
    //output reg out1
);

    //always @(in1) begin
    //    out1 = ?;
    //end

endmodule
